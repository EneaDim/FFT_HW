LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std. all;

ENTITY micro_ROM_odd IS
		PORT(ADDRESS: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
				DATA_OUT_ODD: OUT STD_LOGIC_VECTOR (40 DOWNTO 0));
END micro_ROM_odd;

ARCHITECTURE behaviour OF micro_ROM_odd IS

SIGNAL add: INTEGER RANGE 0 TO 15;
TYPE rom_array_odd IS ARRAY (0 to 15) of STD_LOGIC_VECTOR(40 DOWNTO 0);

CONSTANT ROM: ROM_array_odd:= (
"11001100000000000000000000000000000000000",--RESET
"00001100000011111101110000000011000011110",--S3
"00011100000011111100111111101111000011110",--S6
"00100100000011111101111111011111000011110",--S12
"00110100000011111100010000001111101011110",--S8
"00011100000011111100111111101111000011111",--S15
"01001100000011111100010000000011000011111",--DONE
"00101110101011111110110101011111010111110",--S16
"00010110101011111110110101011111000011110",--S10
"00000110101011111100010000000011000011110",--S1
"00000100000000000000000000000000000000000",--UNDEFINED
"00000100000000000000000000000000000000000",--UNDEFINED
"00000100000000000000000000000000000000000",--UNDEFINED
"00000100000000000000000000000000000000000",--UNDEFINED
"00000100000000000000000000000000000000000",--UNDEFINED
"00000100000000000000000000000000000000000"--UNDEFINED
);
BEGIN 
add <= to_integer(unsigned(ADDRESS));
DATA_OUT_ODD <= ROM(add);
END ARCHITECTURE;