LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std. all;

ENTITY micro_ROM_even IS
		PORT(ADDRESS: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				DATA_OUT_EVEN: OUT STD_LOGIC_VECTOR (40 DOWNTO 0));
END micro_ROM_even;

ARCHITECTURE behaviour OF micro_ROM_even IS

SIGNAL add: INTEGER RANGE 0 TO 15;
TYPE rom_array_even IS ARRAY (0 to 15) of STD_LOGIC_VECTOR(40 DOWNTO 0);

CONSTANT ROM: ROM_array_even:= (
"00001001010111111100010000000011000011110",--S2
"11000000000011111111110000010011000011110",--S4
"00011001010111111100111111101111000011110",--S11
"00100000000011111100011111011111000011110",--S7
"10111000000011111111110000011111101011110",--S13
"00011001010111111100111111101111000011111", --S17
"00110000000011111100010000000011010111110",--S9
"00101000000011111110110101011111010111110",--S14
"00010000000011111110110101011111000011110",--S5
"11001000000011111100010000000011000011110",--IDLE
"00000000000000000000000000000000000000000",--UNDEFINED
"00000000000000000000000000000000000000000",--UNDEFINED
"00000000000000000000000000000000000000000",--UNDEFINED
"00000000000000000000000000000000000000000",--UNDEFINED
"00000000000000000000000000000000000000000",--UNDEFINED
"00000000000000000000000000000000000000000"--UNDEFINED
);
BEGIN 
add <= to_integer(unsigned(ADDRESS));
DATA_OUT_EVEN <= ROM(add);

END ARCHITECTURE;
